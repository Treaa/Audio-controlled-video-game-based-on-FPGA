// nios_cpu.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nios_cpu (
		input  wire        audio_clk_50_clk,                     //           audio_clk_50.clk
		input  wire        audio_io_adc_data,                    //               audio_io.adc_data
		inout  wire        audio_io_adc_clk,                     //                       .adc_clk
		inout  wire        audio_io_bit_stream_clk,              //                       .bit_stream_clk
		output wire        audio_io_dac_data,                    //                       .dac_data
		inout  wire        audio_io_dac_clk,                     //                       .dac_clk
		output wire        audio_io_chip_clk,                    //                       .chip_clk
		output wire        clk_100_clk,                          //                clk_100.clk
		output wire        clk_25_clk,                           //                 clk_25.clk
		input  wire        clk_27_clk,                           //                 clk_27.clk
		input  wire        clk_50_clk,                           //                 clk_50.clk
		output wire        external_i2c_i2c_sclk,                //           external_i2c.i2c_sclk
		inout  wire        external_i2c_i2c_sdat,                //                       .i2c_sdat
		input  wire [3:0]  external_key_key,                     //           external_key.key
		output wire [8:0]  external_led_led,                     //           external_led.led
		output wire [9:0]  external_pio_b_off_export,            //     external_pio_b_off.export
		output wire [9:0]  external_pio_b_on_export,             //      external_pio_b_on.export
		output wire [9:0]  external_pio_g_off_export,            //     external_pio_g_off.export
		output wire [9:0]  external_pio_g_on_export,             //      external_pio_g_on.export
		output wire [18:0] external_pio_pixel_pos_export,        // external_pio_pixel_pos.export
		output wire        external_pio_pos_state_export,        // external_pio_pos_state.export
		output wire [9:0]  external_pio_r_off_export,            //     external_pio_r_off.export
		output wire [9:0]  external_pio_r_on_export,             //      external_pio_r_on.export
		input  wire [2:0]  external_sw_export,                   //            external_sw.export
		input  wire        reset_reset_n,                        //                  reset.reset_n
		output wire [19:0] sram_bridge_out_tcm_address_out,      //        sram_bridge_out.tcm_address_out
		output wire [1:0]  sram_bridge_out_tcm_byteenable_n_out, //                       .tcm_byteenable_n_out
		output wire [0:0]  sram_bridge_out_tcm_read_n_out,       //                       .tcm_read_n_out
		output wire [0:0]  sram_bridge_out_tcm_write_n_out,      //                       .tcm_write_n_out
		inout  wire [15:0] sram_bridge_out_tcm_data_out,         //                       .tcm_data_out
		output wire [0:0]  sram_bridge_out_tcm_chipselect_n_out  //                       .tcm_chipselect_n_out
	);

	wire         pll_100_25_c0_clk;                                           // pll_100_25:c0 -> [audio_process_0:clk, cpu:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:pll_100_25_c0_clk, pio_b_off:clk, pio_b_on:clk, pio_g_off:clk, pio_g_on:clk, pio_pixel_pos:clk, pio_pos_state:clk, pio_r_off:clk, pio_r_on:clk, pio_switch:clk, rst_controller:clk, sram:clk_clk, sram_bridge:clk, sysid_qsys_0:clock, timer:clk]
	wire         sram_tcm_data_outen;                                         // sram:tcm_data_outen -> sram_bridge:tcs_tcm_data_outen
	wire         sram_tcm_request;                                            // sram:tcm_request -> sram_bridge:request
	wire   [1:0] sram_tcm_byteenable_n_out;                                   // sram:tcm_byteenable_n_out -> sram_bridge:tcs_tcm_byteenable_n_out
	wire         sram_tcm_write_n_out;                                        // sram:tcm_write_n_out -> sram_bridge:tcs_tcm_write_n_out
	wire         sram_tcm_read_n_out;                                         // sram:tcm_read_n_out -> sram_bridge:tcs_tcm_read_n_out
	wire         sram_tcm_grant;                                              // sram_bridge:grant -> sram:tcm_grant
	wire         sram_tcm_chipselect_n_out;                                   // sram:tcm_chipselect_n_out -> sram_bridge:tcs_tcm_chipselect_n_out
	wire  [19:0] sram_tcm_address_out;                                        // sram:tcm_address_out -> sram_bridge:tcs_tcm_address_out
	wire  [15:0] sram_tcm_data_out;                                           // sram:tcm_data_out -> sram_bridge:tcs_tcm_data_out
	wire  [15:0] sram_tcm_data_in;                                            // sram_bridge:tcs_tcm_data_in -> sram:tcm_data_in
	wire  [31:0] cpu_data_master_readdata;                                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                 // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [21:0] cpu_data_master_address;                                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                             // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                          // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [21:0] cpu_instruction_master_address;                              // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                 // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                        // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_audio_process_0_avalon_slave_0_chipselect; // mm_interconnect_0:audio_process_0_avalon_slave_0_chipselect -> audio_process_0:chipselect
	wire  [31:0] mm_interconnect_0_audio_process_0_avalon_slave_0_readdata;   // audio_process_0:readdata -> mm_interconnect_0:audio_process_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_audio_process_0_avalon_slave_0_address;    // mm_interconnect_0:audio_process_0_avalon_slave_0_address -> audio_process_0:address
	wire         mm_interconnect_0_audio_process_0_avalon_slave_0_read;       // mm_interconnect_0:audio_process_0_avalon_slave_0_read -> audio_process_0:read
	wire   [3:0] mm_interconnect_0_audio_process_0_avalon_slave_0_byteenable; // mm_interconnect_0:audio_process_0_avalon_slave_0_byteenable -> audio_process_0:byteenable
	wire         mm_interconnect_0_audio_process_0_avalon_slave_0_write;      // mm_interconnect_0:audio_process_0_avalon_slave_0_write -> audio_process_0:write
	wire  [31:0] mm_interconnect_0_audio_process_0_avalon_slave_0_writedata;  // mm_interconnect_0:audio_process_0_avalon_slave_0_writedata -> audio_process_0:writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;              // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;           // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;           // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;               // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                  // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;            // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                 // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;             // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_100_25_pll_slave_readdata;             // pll_100_25:readdata -> mm_interconnect_0:pll_100_25_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_100_25_pll_slave_address;              // mm_interconnect_0:pll_100_25_pll_slave_address -> pll_100_25:address
	wire         mm_interconnect_0_pll_100_25_pll_slave_read;                 // mm_interconnect_0:pll_100_25_pll_slave_read -> pll_100_25:read
	wire         mm_interconnect_0_pll_100_25_pll_slave_write;                // mm_interconnect_0:pll_100_25_pll_slave_write -> pll_100_25:write
	wire  [31:0] mm_interconnect_0_pll_100_25_pll_slave_writedata;            // mm_interconnect_0:pll_100_25_pll_slave_writedata -> pll_100_25:writedata
	wire  [31:0] mm_interconnect_0_pio_switch_s1_readdata;                    // pio_switch:readdata -> mm_interconnect_0:pio_switch_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_switch_s1_address;                     // mm_interconnect_0:pio_switch_s1_address -> pio_switch:address
	wire         mm_interconnect_0_pio_r_on_s1_chipselect;                    // mm_interconnect_0:pio_r_on_s1_chipselect -> pio_r_on:chipselect
	wire  [31:0] mm_interconnect_0_pio_r_on_s1_readdata;                      // pio_r_on:readdata -> mm_interconnect_0:pio_r_on_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_r_on_s1_address;                       // mm_interconnect_0:pio_r_on_s1_address -> pio_r_on:address
	wire         mm_interconnect_0_pio_r_on_s1_write;                         // mm_interconnect_0:pio_r_on_s1_write -> pio_r_on:write_n
	wire  [31:0] mm_interconnect_0_pio_r_on_s1_writedata;                     // mm_interconnect_0:pio_r_on_s1_writedata -> pio_r_on:writedata
	wire         mm_interconnect_0_pio_g_on_s1_chipselect;                    // mm_interconnect_0:pio_g_on_s1_chipselect -> pio_g_on:chipselect
	wire  [31:0] mm_interconnect_0_pio_g_on_s1_readdata;                      // pio_g_on:readdata -> mm_interconnect_0:pio_g_on_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_g_on_s1_address;                       // mm_interconnect_0:pio_g_on_s1_address -> pio_g_on:address
	wire         mm_interconnect_0_pio_g_on_s1_write;                         // mm_interconnect_0:pio_g_on_s1_write -> pio_g_on:write_n
	wire  [31:0] mm_interconnect_0_pio_g_on_s1_writedata;                     // mm_interconnect_0:pio_g_on_s1_writedata -> pio_g_on:writedata
	wire         mm_interconnect_0_pio_b_on_s1_chipselect;                    // mm_interconnect_0:pio_b_on_s1_chipselect -> pio_b_on:chipselect
	wire  [31:0] mm_interconnect_0_pio_b_on_s1_readdata;                      // pio_b_on:readdata -> mm_interconnect_0:pio_b_on_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_b_on_s1_address;                       // mm_interconnect_0:pio_b_on_s1_address -> pio_b_on:address
	wire         mm_interconnect_0_pio_b_on_s1_write;                         // mm_interconnect_0:pio_b_on_s1_write -> pio_b_on:write_n
	wire  [31:0] mm_interconnect_0_pio_b_on_s1_writedata;                     // mm_interconnect_0:pio_b_on_s1_writedata -> pio_b_on:writedata
	wire         mm_interconnect_0_pio_r_off_s1_chipselect;                   // mm_interconnect_0:pio_r_off_s1_chipselect -> pio_r_off:chipselect
	wire  [31:0] mm_interconnect_0_pio_r_off_s1_readdata;                     // pio_r_off:readdata -> mm_interconnect_0:pio_r_off_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_r_off_s1_address;                      // mm_interconnect_0:pio_r_off_s1_address -> pio_r_off:address
	wire         mm_interconnect_0_pio_r_off_s1_write;                        // mm_interconnect_0:pio_r_off_s1_write -> pio_r_off:write_n
	wire  [31:0] mm_interconnect_0_pio_r_off_s1_writedata;                    // mm_interconnect_0:pio_r_off_s1_writedata -> pio_r_off:writedata
	wire         mm_interconnect_0_pio_g_off_s1_chipselect;                   // mm_interconnect_0:pio_g_off_s1_chipselect -> pio_g_off:chipselect
	wire  [31:0] mm_interconnect_0_pio_g_off_s1_readdata;                     // pio_g_off:readdata -> mm_interconnect_0:pio_g_off_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_g_off_s1_address;                      // mm_interconnect_0:pio_g_off_s1_address -> pio_g_off:address
	wire         mm_interconnect_0_pio_g_off_s1_write;                        // mm_interconnect_0:pio_g_off_s1_write -> pio_g_off:write_n
	wire  [31:0] mm_interconnect_0_pio_g_off_s1_writedata;                    // mm_interconnect_0:pio_g_off_s1_writedata -> pio_g_off:writedata
	wire         mm_interconnect_0_pio_b_off_s1_chipselect;                   // mm_interconnect_0:pio_b_off_s1_chipselect -> pio_b_off:chipselect
	wire  [31:0] mm_interconnect_0_pio_b_off_s1_readdata;                     // pio_b_off:readdata -> mm_interconnect_0:pio_b_off_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_b_off_s1_address;                      // mm_interconnect_0:pio_b_off_s1_address -> pio_b_off:address
	wire         mm_interconnect_0_pio_b_off_s1_write;                        // mm_interconnect_0:pio_b_off_s1_write -> pio_b_off:write_n
	wire  [31:0] mm_interconnect_0_pio_b_off_s1_writedata;                    // mm_interconnect_0:pio_b_off_s1_writedata -> pio_b_off:writedata
	wire         mm_interconnect_0_pio_pos_state_s1_chipselect;               // mm_interconnect_0:pio_pos_state_s1_chipselect -> pio_pos_state:chipselect
	wire  [31:0] mm_interconnect_0_pio_pos_state_s1_readdata;                 // pio_pos_state:readdata -> mm_interconnect_0:pio_pos_state_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_pos_state_s1_address;                  // mm_interconnect_0:pio_pos_state_s1_address -> pio_pos_state:address
	wire         mm_interconnect_0_pio_pos_state_s1_write;                    // mm_interconnect_0:pio_pos_state_s1_write -> pio_pos_state:write_n
	wire  [31:0] mm_interconnect_0_pio_pos_state_s1_writedata;                // mm_interconnect_0:pio_pos_state_s1_writedata -> pio_pos_state:writedata
	wire         mm_interconnect_0_pio_pixel_pos_s1_chipselect;               // mm_interconnect_0:pio_pixel_pos_s1_chipselect -> pio_pixel_pos:chipselect
	wire  [31:0] mm_interconnect_0_pio_pixel_pos_s1_readdata;                 // pio_pixel_pos:readdata -> mm_interconnect_0:pio_pixel_pos_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_pixel_pos_s1_address;                  // mm_interconnect_0:pio_pixel_pos_s1_address -> pio_pixel_pos:address
	wire         mm_interconnect_0_pio_pixel_pos_s1_write;                    // mm_interconnect_0:pio_pixel_pos_s1_write -> pio_pixel_pos:write_n
	wire  [31:0] mm_interconnect_0_pio_pixel_pos_s1_writedata;                // mm_interconnect_0:pio_pixel_pos_s1_writedata -> pio_pixel_pos:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                       // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                         // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                          // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                            // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                        // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire  [15:0] mm_interconnect_0_sram_uas_readdata;                         // sram:uas_readdata -> mm_interconnect_0:sram_uas_readdata
	wire         mm_interconnect_0_sram_uas_waitrequest;                      // sram:uas_waitrequest -> mm_interconnect_0:sram_uas_waitrequest
	wire         mm_interconnect_0_sram_uas_debugaccess;                      // mm_interconnect_0:sram_uas_debugaccess -> sram:uas_debugaccess
	wire  [19:0] mm_interconnect_0_sram_uas_address;                          // mm_interconnect_0:sram_uas_address -> sram:uas_address
	wire         mm_interconnect_0_sram_uas_read;                             // mm_interconnect_0:sram_uas_read -> sram:uas_read
	wire   [1:0] mm_interconnect_0_sram_uas_byteenable;                       // mm_interconnect_0:sram_uas_byteenable -> sram:uas_byteenable
	wire         mm_interconnect_0_sram_uas_readdatavalid;                    // sram:uas_readdatavalid -> mm_interconnect_0:sram_uas_readdatavalid
	wire         mm_interconnect_0_sram_uas_lock;                             // mm_interconnect_0:sram_uas_lock -> sram:uas_lock
	wire         mm_interconnect_0_sram_uas_write;                            // mm_interconnect_0:sram_uas_write -> sram:uas_write
	wire  [15:0] mm_interconnect_0_sram_uas_writedata;                        // mm_interconnect_0:sram_uas_writedata -> sram:uas_writedata
	wire   [1:0] mm_interconnect_0_sram_uas_burstcount;                       // mm_interconnect_0:sram_uas_burstcount -> sram:uas_burstcount
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // timer:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                                 // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [audio_process_0:reset_n, cpu:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, pio_b_off:reset_n, pio_b_on:reset_n, pio_g_off:reset_n, pio_g_on:reset_n, pio_pixel_pos:reset_n, pio_pos_state:reset_n, pio_r_off:reset_n, pio_r_on:reset_n, pio_switch:reset_n, rst_translator:in_reset, sram:reset_reset, sram_bridge:reset, sysid_qsys_0:reset_n, timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [mm_interconnect_0:pll_100_25_inclk_interface_reset_reset_bridge_in_reset_reset, pll_100_25:reset]

	audio_proc_avalon_mm audio_process_0 (
		.address     (mm_interconnect_0_audio_process_0_avalon_slave_0_address),    //    avalon_slave_0.address
		.writedata   (mm_interconnect_0_audio_process_0_avalon_slave_0_writedata),  //                  .writedata
		.byteenable  (mm_interconnect_0_audio_process_0_avalon_slave_0_byteenable), //                  .byteenable
		.write       (mm_interconnect_0_audio_process_0_avalon_slave_0_write),      //                  .write
		.read        (mm_interconnect_0_audio_process_0_avalon_slave_0_read),       //                  .read
		.chipselect  (mm_interconnect_0_audio_process_0_avalon_slave_0_chipselect), //                  .chipselect
		.readdata    (mm_interconnect_0_audio_process_0_avalon_slave_0_readdata),   //                  .readdata
		.AUD_ADCDAT  (audio_io_adc_data),                                           // external_audio_io.adc_data
		.AUD_ADCLRCK (audio_io_adc_clk),                                            //                  .adc_clk
		.AUD_BCLK    (audio_io_bit_stream_clk),                                     //                  .bit_stream_clk
		.AUD_DACDAT  (audio_io_dac_data),                                           //                  .dac_data
		.AUD_DACLRCK (audio_io_dac_clk),                                            //                  .dac_clk
		.AUD_XCK     (audio_io_chip_clk),                                           //                  .chip_clk
		.clk         (pll_100_25_c0_clk),                                           //               clk.clk
		.CLOCK_27    (clk_27_clk),                                                  //            clk_27.clk
		.CLOCK_50    (audio_clk_50_clk),                                            //            clk_50.clk
		.LEDG        (external_led_led),                                            //      external_led.led
		.KEY         (external_key_key),                                            //      external_key.key
		.reset_n     (~rst_controller_reset_out_reset),                             //           reset_n.reset_n
		.I2C_SCLK    (external_i2c_i2c_sclk),                                       //      external_I2C.i2c_sclk
		.I2C_SDAT    (external_i2c_i2c_sdat)                                        //                  .i2c_sdat
	);

	nios_cpu_cpu cpu (
		.clk                                 (pll_100_25_c0_clk),                                 //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	nios_cpu_jtag_uart_0 jtag_uart_0 (
		.clk            (pll_100_25_c0_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	nios_cpu_pio_b_off pio_b_off (
		.clk        (pll_100_25_c0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_b_off_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_b_off_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_b_off_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_b_off_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_b_off_s1_readdata),   //                    .readdata
		.out_port   (external_pio_b_off_export)                  // external_connection.export
	);

	nios_cpu_pio_b_off pio_b_on (
		.clk        (pll_100_25_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_pio_b_on_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_b_on_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_b_on_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_b_on_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_b_on_s1_readdata),   //                    .readdata
		.out_port   (external_pio_b_on_export)                  // external_connection.export
	);

	nios_cpu_pio_b_off pio_g_off (
		.clk        (pll_100_25_c0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_g_off_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_g_off_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_g_off_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_g_off_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_g_off_s1_readdata),   //                    .readdata
		.out_port   (external_pio_g_off_export)                  // external_connection.export
	);

	nios_cpu_pio_b_off pio_g_on (
		.clk        (pll_100_25_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_pio_g_on_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_g_on_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_g_on_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_g_on_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_g_on_s1_readdata),   //                    .readdata
		.out_port   (external_pio_g_on_export)                  // external_connection.export
	);

	nios_cpu_pio_pixel_pos pio_pixel_pos (
		.clk        (pll_100_25_c0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_pixel_pos_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_pixel_pos_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_pixel_pos_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_pixel_pos_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_pixel_pos_s1_readdata),   //                    .readdata
		.out_port   (external_pio_pixel_pos_export)                  // external_connection.export
	);

	nios_cpu_pio_pos_state pio_pos_state (
		.clk        (pll_100_25_c0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_pos_state_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_pos_state_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_pos_state_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_pos_state_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_pos_state_s1_readdata),   //                    .readdata
		.out_port   (external_pio_pos_state_export)                  // external_connection.export
	);

	nios_cpu_pio_b_off pio_r_off (
		.clk        (pll_100_25_c0_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_r_off_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_r_off_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_r_off_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_r_off_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_r_off_s1_readdata),   //                    .readdata
		.out_port   (external_pio_r_off_export)                  // external_connection.export
	);

	nios_cpu_pio_b_off pio_r_on (
		.clk        (pll_100_25_c0_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_pio_r_on_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_r_on_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_r_on_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_r_on_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_r_on_s1_readdata),   //                    .readdata
		.out_port   (external_pio_r_on_export)                  // external_connection.export
	);

	nios_cpu_pio_switch pio_switch (
		.clk      (pll_100_25_c0_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pio_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_switch_s1_readdata), //                    .readdata
		.in_port  (external_sw_export)                        // external_connection.export
	);

	nios_cpu_pll_100_25 pll_100_25 (
		.clk                (clk_50_clk),                                       //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),               // inclk_interface_reset.reset
		.read               (mm_interconnect_0_pll_100_25_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_pll_100_25_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_pll_100_25_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_pll_100_25_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_pll_100_25_pll_slave_writedata), //                      .writedata
		.c0                 (pll_100_25_c0_clk),                                //                    c0.clk
		.c1                 (clk_25_clk),                                       //                    c1.clk
		.c2                 (clk_100_clk),                                      //                    c2.clk
		.scandone           (),                                                 //           (terminated)
		.scandataout        (),                                                 //           (terminated)
		.areset             (1'b0),                                             //           (terminated)
		.locked             (),                                                 //           (terminated)
		.phasedone          (),                                                 //           (terminated)
		.phasecounterselect (4'b0000),                                          //           (terminated)
		.phaseupdown        (1'b0),                                             //           (terminated)
		.phasestep          (1'b0),                                             //           (terminated)
		.scanclk            (1'b0),                                             //           (terminated)
		.scanclkena         (1'b0),                                             //           (terminated)
		.scandata           (1'b0),                                             //           (terminated)
		.configupdate       (1'b0)                                              //           (terminated)
	);

	nios_cpu_sram #(
		.TCM_ADDRESS_W                  (20),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (20),
		.TCM_WRITE_WAIT                 (10),
		.TCM_SETUP_WAIT                 (5),
		.TCM_DATA_HOLD                  (10),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) sram (
		.clk_clk              (pll_100_25_c0_clk),                        //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),           // reset.reset
		.uas_address          (mm_interconnect_0_sram_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_sram_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_sram_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_sram_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_sram_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_sram_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_sram_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_sram_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_sram_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_sram_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_sram_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (sram_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (sram_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (sram_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (sram_tcm_request),                         //      .request
		.tcm_grant            (sram_tcm_grant),                           //      .grant
		.tcm_address_out      (sram_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out (sram_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out         (sram_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (sram_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (sram_tcm_data_in)                          //      .data_in
	);

	nios_cpu_sram_bridge sram_bridge (
		.clk                      (pll_100_25_c0_clk),                    //   clk.clk
		.reset                    (rst_controller_reset_out_reset),       // reset.reset
		.request                  (sram_tcm_request),                     //   tcs.request
		.grant                    (sram_tcm_grant),                       //      .grant
		.tcs_tcm_address_out      (sram_tcm_address_out),                 //      .address_out
		.tcs_tcm_byteenable_n_out (sram_tcm_byteenable_n_out),            //      .byteenable_n_out
		.tcs_tcm_read_n_out       (sram_tcm_read_n_out),                  //      .read_n_out
		.tcs_tcm_write_n_out      (sram_tcm_write_n_out),                 //      .write_n_out
		.tcs_tcm_data_out         (sram_tcm_data_out),                    //      .data_out
		.tcs_tcm_data_outen       (sram_tcm_data_outen),                  //      .data_outen
		.tcs_tcm_data_in          (sram_tcm_data_in),                     //      .data_in
		.tcs_tcm_chipselect_n_out (sram_tcm_chipselect_n_out),            //      .chipselect_n_out
		.tcm_address_out          (sram_bridge_out_tcm_address_out),      //   out.tcm_address_out
		.tcm_byteenable_n_out     (sram_bridge_out_tcm_byteenable_n_out), //      .tcm_byteenable_n_out
		.tcm_read_n_out           (sram_bridge_out_tcm_read_n_out),       //      .tcm_read_n_out
		.tcm_write_n_out          (sram_bridge_out_tcm_write_n_out),      //      .tcm_write_n_out
		.tcm_data_out             (sram_bridge_out_tcm_data_out),         //      .tcm_data_out
		.tcm_chipselect_n_out     (sram_bridge_out_tcm_chipselect_n_out)  //      .tcm_chipselect_n_out
	);

	nios_cpu_sysid_qsys_0 sysid_qsys_0 (
		.clock    (pll_100_25_c0_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_cpu_timer timer (
		.clk        (pll_100_25_c0_clk),                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	nios_cpu_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                (clk_50_clk),                                                  //                                              clk_0_clk.clk
		.pll_100_25_c0_clk                                            (pll_100_25_c0_clk),                                           //                                          pll_100_25_c0.clk
		.cpu_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                              //                        cpu_reset_reset_bridge_in_reset.reset
		.pll_100_25_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // pll_100_25_inclk_interface_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                      (cpu_data_master_address),                                     //                                        cpu_data_master.address
		.cpu_data_master_waitrequest                                  (cpu_data_master_waitrequest),                                 //                                                       .waitrequest
		.cpu_data_master_byteenable                                   (cpu_data_master_byteenable),                                  //                                                       .byteenable
		.cpu_data_master_read                                         (cpu_data_master_read),                                        //                                                       .read
		.cpu_data_master_readdata                                     (cpu_data_master_readdata),                                    //                                                       .readdata
		.cpu_data_master_write                                        (cpu_data_master_write),                                       //                                                       .write
		.cpu_data_master_writedata                                    (cpu_data_master_writedata),                                   //                                                       .writedata
		.cpu_data_master_debugaccess                                  (cpu_data_master_debugaccess),                                 //                                                       .debugaccess
		.cpu_instruction_master_address                               (cpu_instruction_master_address),                              //                                 cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                           (cpu_instruction_master_waitrequest),                          //                                                       .waitrequest
		.cpu_instruction_master_read                                  (cpu_instruction_master_read),                                 //                                                       .read
		.cpu_instruction_master_readdata                              (cpu_instruction_master_readdata),                             //                                                       .readdata
		.cpu_instruction_master_readdatavalid                         (cpu_instruction_master_readdatavalid),                        //                                                       .readdatavalid
		.audio_process_0_avalon_slave_0_address                       (mm_interconnect_0_audio_process_0_avalon_slave_0_address),    //                         audio_process_0_avalon_slave_0.address
		.audio_process_0_avalon_slave_0_write                         (mm_interconnect_0_audio_process_0_avalon_slave_0_write),      //                                                       .write
		.audio_process_0_avalon_slave_0_read                          (mm_interconnect_0_audio_process_0_avalon_slave_0_read),       //                                                       .read
		.audio_process_0_avalon_slave_0_readdata                      (mm_interconnect_0_audio_process_0_avalon_slave_0_readdata),   //                                                       .readdata
		.audio_process_0_avalon_slave_0_writedata                     (mm_interconnect_0_audio_process_0_avalon_slave_0_writedata),  //                                                       .writedata
		.audio_process_0_avalon_slave_0_byteenable                    (mm_interconnect_0_audio_process_0_avalon_slave_0_byteenable), //                                                       .byteenable
		.audio_process_0_avalon_slave_0_chipselect                    (mm_interconnect_0_audio_process_0_avalon_slave_0_chipselect), //                                                       .chipselect
		.cpu_debug_mem_slave_address                                  (mm_interconnect_0_cpu_debug_mem_slave_address),               //                                    cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                    (mm_interconnect_0_cpu_debug_mem_slave_write),                 //                                                       .write
		.cpu_debug_mem_slave_read                                     (mm_interconnect_0_cpu_debug_mem_slave_read),                  //                                                       .read
		.cpu_debug_mem_slave_readdata                                 (mm_interconnect_0_cpu_debug_mem_slave_readdata),              //                                                       .readdata
		.cpu_debug_mem_slave_writedata                                (mm_interconnect_0_cpu_debug_mem_slave_writedata),             //                                                       .writedata
		.cpu_debug_mem_slave_byteenable                               (mm_interconnect_0_cpu_debug_mem_slave_byteenable),            //                                                       .byteenable
		.cpu_debug_mem_slave_waitrequest                              (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),           //                                                       .waitrequest
		.cpu_debug_mem_slave_debugaccess                              (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),           //                                                       .debugaccess
		.jtag_uart_0_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                          jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                                       .write
		.jtag_uart_0_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                                       .read
		.jtag_uart_0_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                                       .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                                       .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                                       .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                                       .chipselect
		.pio_b_off_s1_address                                         (mm_interconnect_0_pio_b_off_s1_address),                      //                                           pio_b_off_s1.address
		.pio_b_off_s1_write                                           (mm_interconnect_0_pio_b_off_s1_write),                        //                                                       .write
		.pio_b_off_s1_readdata                                        (mm_interconnect_0_pio_b_off_s1_readdata),                     //                                                       .readdata
		.pio_b_off_s1_writedata                                       (mm_interconnect_0_pio_b_off_s1_writedata),                    //                                                       .writedata
		.pio_b_off_s1_chipselect                                      (mm_interconnect_0_pio_b_off_s1_chipselect),                   //                                                       .chipselect
		.pio_b_on_s1_address                                          (mm_interconnect_0_pio_b_on_s1_address),                       //                                            pio_b_on_s1.address
		.pio_b_on_s1_write                                            (mm_interconnect_0_pio_b_on_s1_write),                         //                                                       .write
		.pio_b_on_s1_readdata                                         (mm_interconnect_0_pio_b_on_s1_readdata),                      //                                                       .readdata
		.pio_b_on_s1_writedata                                        (mm_interconnect_0_pio_b_on_s1_writedata),                     //                                                       .writedata
		.pio_b_on_s1_chipselect                                       (mm_interconnect_0_pio_b_on_s1_chipselect),                    //                                                       .chipselect
		.pio_g_off_s1_address                                         (mm_interconnect_0_pio_g_off_s1_address),                      //                                           pio_g_off_s1.address
		.pio_g_off_s1_write                                           (mm_interconnect_0_pio_g_off_s1_write),                        //                                                       .write
		.pio_g_off_s1_readdata                                        (mm_interconnect_0_pio_g_off_s1_readdata),                     //                                                       .readdata
		.pio_g_off_s1_writedata                                       (mm_interconnect_0_pio_g_off_s1_writedata),                    //                                                       .writedata
		.pio_g_off_s1_chipselect                                      (mm_interconnect_0_pio_g_off_s1_chipselect),                   //                                                       .chipselect
		.pio_g_on_s1_address                                          (mm_interconnect_0_pio_g_on_s1_address),                       //                                            pio_g_on_s1.address
		.pio_g_on_s1_write                                            (mm_interconnect_0_pio_g_on_s1_write),                         //                                                       .write
		.pio_g_on_s1_readdata                                         (mm_interconnect_0_pio_g_on_s1_readdata),                      //                                                       .readdata
		.pio_g_on_s1_writedata                                        (mm_interconnect_0_pio_g_on_s1_writedata),                     //                                                       .writedata
		.pio_g_on_s1_chipselect                                       (mm_interconnect_0_pio_g_on_s1_chipselect),                    //                                                       .chipselect
		.pio_pixel_pos_s1_address                                     (mm_interconnect_0_pio_pixel_pos_s1_address),                  //                                       pio_pixel_pos_s1.address
		.pio_pixel_pos_s1_write                                       (mm_interconnect_0_pio_pixel_pos_s1_write),                    //                                                       .write
		.pio_pixel_pos_s1_readdata                                    (mm_interconnect_0_pio_pixel_pos_s1_readdata),                 //                                                       .readdata
		.pio_pixel_pos_s1_writedata                                   (mm_interconnect_0_pio_pixel_pos_s1_writedata),                //                                                       .writedata
		.pio_pixel_pos_s1_chipselect                                  (mm_interconnect_0_pio_pixel_pos_s1_chipselect),               //                                                       .chipselect
		.pio_pos_state_s1_address                                     (mm_interconnect_0_pio_pos_state_s1_address),                  //                                       pio_pos_state_s1.address
		.pio_pos_state_s1_write                                       (mm_interconnect_0_pio_pos_state_s1_write),                    //                                                       .write
		.pio_pos_state_s1_readdata                                    (mm_interconnect_0_pio_pos_state_s1_readdata),                 //                                                       .readdata
		.pio_pos_state_s1_writedata                                   (mm_interconnect_0_pio_pos_state_s1_writedata),                //                                                       .writedata
		.pio_pos_state_s1_chipselect                                  (mm_interconnect_0_pio_pos_state_s1_chipselect),               //                                                       .chipselect
		.pio_r_off_s1_address                                         (mm_interconnect_0_pio_r_off_s1_address),                      //                                           pio_r_off_s1.address
		.pio_r_off_s1_write                                           (mm_interconnect_0_pio_r_off_s1_write),                        //                                                       .write
		.pio_r_off_s1_readdata                                        (mm_interconnect_0_pio_r_off_s1_readdata),                     //                                                       .readdata
		.pio_r_off_s1_writedata                                       (mm_interconnect_0_pio_r_off_s1_writedata),                    //                                                       .writedata
		.pio_r_off_s1_chipselect                                      (mm_interconnect_0_pio_r_off_s1_chipselect),                   //                                                       .chipselect
		.pio_r_on_s1_address                                          (mm_interconnect_0_pio_r_on_s1_address),                       //                                            pio_r_on_s1.address
		.pio_r_on_s1_write                                            (mm_interconnect_0_pio_r_on_s1_write),                         //                                                       .write
		.pio_r_on_s1_readdata                                         (mm_interconnect_0_pio_r_on_s1_readdata),                      //                                                       .readdata
		.pio_r_on_s1_writedata                                        (mm_interconnect_0_pio_r_on_s1_writedata),                     //                                                       .writedata
		.pio_r_on_s1_chipselect                                       (mm_interconnect_0_pio_r_on_s1_chipselect),                    //                                                       .chipselect
		.pio_switch_s1_address                                        (mm_interconnect_0_pio_switch_s1_address),                     //                                          pio_switch_s1.address
		.pio_switch_s1_readdata                                       (mm_interconnect_0_pio_switch_s1_readdata),                    //                                                       .readdata
		.pll_100_25_pll_slave_address                                 (mm_interconnect_0_pll_100_25_pll_slave_address),              //                                   pll_100_25_pll_slave.address
		.pll_100_25_pll_slave_write                                   (mm_interconnect_0_pll_100_25_pll_slave_write),                //                                                       .write
		.pll_100_25_pll_slave_read                                    (mm_interconnect_0_pll_100_25_pll_slave_read),                 //                                                       .read
		.pll_100_25_pll_slave_readdata                                (mm_interconnect_0_pll_100_25_pll_slave_readdata),             //                                                       .readdata
		.pll_100_25_pll_slave_writedata                               (mm_interconnect_0_pll_100_25_pll_slave_writedata),            //                                                       .writedata
		.sram_uas_address                                             (mm_interconnect_0_sram_uas_address),                          //                                               sram_uas.address
		.sram_uas_write                                               (mm_interconnect_0_sram_uas_write),                            //                                                       .write
		.sram_uas_read                                                (mm_interconnect_0_sram_uas_read),                             //                                                       .read
		.sram_uas_readdata                                            (mm_interconnect_0_sram_uas_readdata),                         //                                                       .readdata
		.sram_uas_writedata                                           (mm_interconnect_0_sram_uas_writedata),                        //                                                       .writedata
		.sram_uas_burstcount                                          (mm_interconnect_0_sram_uas_burstcount),                       //                                                       .burstcount
		.sram_uas_byteenable                                          (mm_interconnect_0_sram_uas_byteenable),                       //                                                       .byteenable
		.sram_uas_readdatavalid                                       (mm_interconnect_0_sram_uas_readdatavalid),                    //                                                       .readdatavalid
		.sram_uas_waitrequest                                         (mm_interconnect_0_sram_uas_waitrequest),                      //                                                       .waitrequest
		.sram_uas_lock                                                (mm_interconnect_0_sram_uas_lock),                             //                                                       .lock
		.sram_uas_debugaccess                                         (mm_interconnect_0_sram_uas_debugaccess),                      //                                                       .debugaccess
		.sysid_qsys_0_control_slave_address                           (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //                             sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                          (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),       //                                                       .readdata
		.timer_s1_address                                             (mm_interconnect_0_timer_s1_address),                          //                                               timer_s1.address
		.timer_s1_write                                               (mm_interconnect_0_timer_s1_write),                            //                                                       .write
		.timer_s1_readdata                                            (mm_interconnect_0_timer_s1_readdata),                         //                                                       .readdata
		.timer_s1_writedata                                           (mm_interconnect_0_timer_s1_writedata),                        //                                                       .writedata
		.timer_s1_chipselect                                          (mm_interconnect_0_timer_s1_chipselect)                        //                                                       .chipselect
	);

	nios_cpu_irq_mapper irq_mapper (
		.clk           (pll_100_25_c0_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_100_25_c0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_50_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
