// Infer ROM storage for a hanning window
module hanningrom (
    input      [9:0]  iAddress,
    output reg [15:0] oHanning
);

always @ (iAddress)
begin
    case (iAddress)
        10'h00: oHanning = 16'h000;
        10'h01: oHanning = 16'h000;
        10'h02: oHanning = 16'h000;
        10'h03: oHanning = 16'h001;
        10'h04: oHanning = 16'h001;
        10'h05: oHanning = 16'h002;
        10'h06: oHanning = 16'h003;
        10'h07: oHanning = 16'h004;
        10'h08: oHanning = 16'h006;
        10'h09: oHanning = 16'h007;
        10'h0a: oHanning = 16'h009;
        10'h0b: oHanning = 16'h00b;
        10'h0c: oHanning = 16'h00c;
        10'h0d: oHanning = 16'h00f;
        10'h0e: oHanning = 16'h011;
        10'h0f: oHanning = 16'h013;
        10'h10: oHanning = 16'h016;
        10'h11: oHanning = 16'h018;
        10'h12: oHanning = 16'h01b;
        10'h13: oHanning = 16'h01e;
        10'h14: oHanning = 16'h021;
        10'h15: oHanning = 16'h025;
        10'h16: oHanning = 16'h028;
        10'h17: oHanning = 16'h02c;
        10'h18: oHanning = 16'h030;
        10'h19: oHanning = 16'h033;
        10'h1a: oHanning = 16'h037;
        10'h1b: oHanning = 16'h03c;
        10'h1c: oHanning = 16'h040;
        10'h1d: oHanning = 16'h045;
        10'h1e: oHanning = 16'h049;
        10'h1f: oHanning = 16'h04e;
        10'h20: oHanning = 16'h053;
        10'h21: oHanning = 16'h058;
        10'h22: oHanning = 16'h05d;
        10'h23: oHanning = 16'h063;
        10'h24: oHanning = 16'h068;
        10'h25: oHanning = 16'h06e;
        10'h26: oHanning = 16'h074;
        10'h27: oHanning = 16'h07a;
        10'h28: oHanning = 16'h080;
        10'h29: oHanning = 16'h087;
        10'h2a: oHanning = 16'h08d;
        10'h2b: oHanning = 16'h094;
        10'h2c: oHanning = 16'h09a;
        10'h2d: oHanning = 16'h0a1;
        10'h2e: oHanning = 16'h0a8;
        10'h2f: oHanning = 16'h0b0;
        10'h30: oHanning = 16'h0b7;
        10'h31: oHanning = 16'h0be;
        10'h32: oHanning = 16'h0c6;
        10'h33: oHanning = 16'h0ce;
        10'h34: oHanning = 16'h0d6;
        10'h35: oHanning = 16'h0de;
        10'h36: oHanning = 16'h0e6;
        10'h37: oHanning = 16'h0ee;
        10'h38: oHanning = 16'h0f7;
        10'h39: oHanning = 16'h100;
        10'h3a: oHanning = 16'h108;
        10'h3b: oHanning = 16'h111;
        10'h3c: oHanning = 16'h11b;
        10'h3d: oHanning = 16'h124;
        10'h3e: oHanning = 16'h12d;
        10'h3f: oHanning = 16'h137;
        10'h40: oHanning = 16'h140;
        10'h41: oHanning = 16'h14a;
        10'h42: oHanning = 16'h154;
        10'h43: oHanning = 16'h15e;
        10'h44: oHanning = 16'h168;
        10'h45: oHanning = 16'h173;
        10'h46: oHanning = 16'h17d;
        10'h47: oHanning = 16'h188;
        10'h48: oHanning = 16'h193;
        10'h49: oHanning = 16'h19e;
        10'h4a: oHanning = 16'h1a9;
        10'h4b: oHanning = 16'h1b4;
        10'h4c: oHanning = 16'h1bf;
        10'h4d: oHanning = 16'h1cb;
        10'h4e: oHanning = 16'h1d6;
        10'h4f: oHanning = 16'h1e2;
        10'h50: oHanning = 16'h1ee;
        10'h51: oHanning = 16'h1fa;
        10'h52: oHanning = 16'h206;
        10'h53: oHanning = 16'h213;
        10'h54: oHanning = 16'h21f;
        10'h55: oHanning = 16'h22c;
        10'h56: oHanning = 16'h238;
        10'h57: oHanning = 16'h245;
        10'h58: oHanning = 16'h252;
        10'h59: oHanning = 16'h25f;
        10'h5a: oHanning = 16'h26c;
        10'h5b: oHanning = 16'h27a;
        10'h5c: oHanning = 16'h287;
        10'h5d: oHanning = 16'h295;
        10'h5e: oHanning = 16'h2a3;
        10'h5f: oHanning = 16'h2b0;
        10'h60: oHanning = 16'h2be;
        10'h61: oHanning = 16'h2cd;
        10'h62: oHanning = 16'h2db;
        10'h63: oHanning = 16'h2e9;
        10'h64: oHanning = 16'h2f8;
        10'h65: oHanning = 16'h306;
        10'h66: oHanning = 16'h315;
        10'h67: oHanning = 16'h324;
        10'h68: oHanning = 16'h333;
        10'h69: oHanning = 16'h342;
        10'h6a: oHanning = 16'h351;
        10'h6b: oHanning = 16'h361;
        10'h6c: oHanning = 16'h370;
        10'h6d: oHanning = 16'h380;
        10'h6e: oHanning = 16'h390;
        10'h6f: oHanning = 16'h3a0;
        10'h70: oHanning = 16'h3af;
        10'h71: oHanning = 16'h3c0;
        10'h72: oHanning = 16'h3d0;
        10'h73: oHanning = 16'h3e0;
        10'h74: oHanning = 16'h3f1;
        10'h75: oHanning = 16'h401;
        10'h76: oHanning = 16'h412;
        10'h77: oHanning = 16'h423;
        10'h78: oHanning = 16'h433;
        10'h79: oHanning = 16'h445;
        10'h7a: oHanning = 16'h456;
        10'h7b: oHanning = 16'h467;
        10'h7c: oHanning = 16'h478;
        10'h7d: oHanning = 16'h48a;
        10'h7e: oHanning = 16'h49b;
        10'h7f: oHanning = 16'h4ad;
        10'h80: oHanning = 16'h4bf;
        10'h81: oHanning = 16'h4d1;
        10'h82: oHanning = 16'h4e3;
        10'h83: oHanning = 16'h4f5;
        10'h84: oHanning = 16'h507;
        10'h85: oHanning = 16'h519;
        10'h86: oHanning = 16'h52c;
        10'h87: oHanning = 16'h53e;
        10'h88: oHanning = 16'h551;
        10'h89: oHanning = 16'h564;
        10'h8a: oHanning = 16'h577;
        10'h8b: oHanning = 16'h58a;
        10'h8c: oHanning = 16'h59d;
        10'h8d: oHanning = 16'h5b0;
        10'h8e: oHanning = 16'h5c3;
        10'h8f: oHanning = 16'h5d6;
        10'h90: oHanning = 16'h5ea;
        10'h91: oHanning = 16'h5fd;
        10'h92: oHanning = 16'h611;
        10'h93: oHanning = 16'h625;
        10'h94: oHanning = 16'h638;
        10'h95: oHanning = 16'h64c;
        10'h96: oHanning = 16'h660;
        10'h97: oHanning = 16'h675;
        10'h98: oHanning = 16'h689;
        10'h99: oHanning = 16'h69d;
        10'h9a: oHanning = 16'h6b1;
        10'h9b: oHanning = 16'h6c6;
        10'h9c: oHanning = 16'h6da;
        10'h9d: oHanning = 16'h6ef;
        10'h9e: oHanning = 16'h704;
        10'h9f: oHanning = 16'h719;
        10'ha0: oHanning = 16'h72e;
        10'ha1: oHanning = 16'h743;
        10'ha2: oHanning = 16'h758;
        10'ha3: oHanning = 16'h76d;
        10'ha4: oHanning = 16'h782;
        10'ha5: oHanning = 16'h797;
        10'ha6: oHanning = 16'h7ad;
        10'ha7: oHanning = 16'h7c2;
        10'ha8: oHanning = 16'h7d8;
        10'ha9: oHanning = 16'h7ed;
        10'haa: oHanning = 16'h803;
        10'hab: oHanning = 16'h819;
        10'hac: oHanning = 16'h82f;
        10'had: oHanning = 16'h845;
        10'hae: oHanning = 16'h85b;
        10'haf: oHanning = 16'h871;
        10'hb0: oHanning = 16'h887;
        10'hb1: oHanning = 16'h89d;
        10'hb2: oHanning = 16'h8b4;
        10'hb3: oHanning = 16'h8ca;
        10'hb4: oHanning = 16'h8e0;
        10'hb5: oHanning = 16'h8f7;
        10'hb6: oHanning = 16'h90e;
        10'hb7: oHanning = 16'h924;
        10'hb8: oHanning = 16'h93b;
        10'hb9: oHanning = 16'h952;
        10'hba: oHanning = 16'h969;
        10'hbb: oHanning = 16'h97f;
        10'hbc: oHanning = 16'h996;
        10'hbd: oHanning = 16'h9ad;
        10'hbe: oHanning = 16'h9c5;
        10'hbf: oHanning = 16'h9dc;
        10'hc0: oHanning = 16'h9f3;
        10'hc1: oHanning = 16'ha0a;
        10'hc2: oHanning = 16'ha21;
        10'hc3: oHanning = 16'ha39;
        10'hc4: oHanning = 16'ha50;
        10'hc5: oHanning = 16'ha68;
        10'hc6: oHanning = 16'ha7f;
        10'hc7: oHanning = 16'ha97;
        10'hc8: oHanning = 16'haaf;
        10'hc9: oHanning = 16'hac6;
        10'hca: oHanning = 16'hade;
        10'hcb: oHanning = 16'haf6;
        10'hcc: oHanning = 16'hb0e;
        10'hcd: oHanning = 16'hb26;
        10'hce: oHanning = 16'hb3e;
        10'hcf: oHanning = 16'hb56;
        10'hd0: oHanning = 16'hb6e;
        10'hd1: oHanning = 16'hb86;
        10'hd2: oHanning = 16'hb9e;
        10'hd3: oHanning = 16'hbb6;
        10'hd4: oHanning = 16'hbce;
        10'hd5: oHanning = 16'hbe6;
        10'hd6: oHanning = 16'hbff;
        10'hd7: oHanning = 16'hc17;
        10'hd8: oHanning = 16'hc2f;
        10'hd9: oHanning = 16'hc48;
        10'hda: oHanning = 16'hc60;
        10'hdb: oHanning = 16'hc79;
        10'hdc: oHanning = 16'hc91;
        10'hdd: oHanning = 16'hcaa;
        10'hde: oHanning = 16'hcc2;
        10'hdf: oHanning = 16'hcdb;
        10'he0: oHanning = 16'hcf4;
        10'he1: oHanning = 16'hd0c;
        10'he2: oHanning = 16'hd25;
        10'he3: oHanning = 16'hd3e;
        10'he4: oHanning = 16'hd56;
        10'he5: oHanning = 16'hd6f;
        10'he6: oHanning = 16'hd88;
        10'he7: oHanning = 16'hda1;
        10'he8: oHanning = 16'hdba;
        10'he9: oHanning = 16'hdd3;
        10'hea: oHanning = 16'hdeb;
        10'heb: oHanning = 16'he04;
        10'hec: oHanning = 16'he1d;
        10'hed: oHanning = 16'he36;
        10'hee: oHanning = 16'he4f;
        10'hef: oHanning = 16'he68;
        10'hf0: oHanning = 16'he81;
        10'hf1: oHanning = 16'he9a;
        10'hf2: oHanning = 16'heb3;
        10'hf3: oHanning = 16'hecc;
        10'hf4: oHanning = 16'hee5;
        10'hf5: oHanning = 16'hefe;
        10'hf6: oHanning = 16'hf17;
        10'hf7: oHanning = 16'hf30;
        10'hf8: oHanning = 16'hf4a;
        10'hf9: oHanning = 16'hf63;
        10'hfa: oHanning = 16'hf7c;
        10'hfb: oHanning = 16'hf95;
        10'hfc: oHanning = 16'hfae;
        10'hfd: oHanning = 16'hfc7;
        10'hfe: oHanning = 16'hfe0;
        10'hff: oHanning = 16'hff9;
        10'h100: oHanning = 16'h1012;
        10'h101: oHanning = 16'h102b;
        10'h102: oHanning = 16'h1045;
        10'h103: oHanning = 16'h105e;
        10'h104: oHanning = 16'h1077;
        10'h105: oHanning = 16'h1090;
        10'h106: oHanning = 16'h10a9;
        10'h107: oHanning = 16'h10c2;
        10'h108: oHanning = 16'h10db;
        10'h109: oHanning = 16'h10f4;
        10'h10a: oHanning = 16'h110d;
        10'h10b: oHanning = 16'h1126;
        10'h10c: oHanning = 16'h113f;
        10'h10d: oHanning = 16'h1158;
        10'h10e: oHanning = 16'h1171;
        10'h10f: oHanning = 16'h118a;
        10'h110: oHanning = 16'h11a3;
        10'h111: oHanning = 16'h11bc;
        10'h112: oHanning = 16'h11d5;
        10'h113: oHanning = 16'h11ee;
        10'h114: oHanning = 16'h1207;
        10'h115: oHanning = 16'h1220;
        10'h116: oHanning = 16'h1239;
        10'h117: oHanning = 16'h1252;
        10'h118: oHanning = 16'h126b;
        10'h119: oHanning = 16'h1283;
        10'h11a: oHanning = 16'h129c;
        10'h11b: oHanning = 16'h12b5;
        10'h11c: oHanning = 16'h12ce;
        10'h11d: oHanning = 16'h12e6;
        10'h11e: oHanning = 16'h12ff;
        10'h11f: oHanning = 16'h1318;
        10'h120: oHanning = 16'h1330;
        10'h121: oHanning = 16'h1349;
        10'h122: oHanning = 16'h1361;
        10'h123: oHanning = 16'h137a;
        10'h124: oHanning = 16'h1392;
        10'h125: oHanning = 16'h13ab;
        10'h126: oHanning = 16'h13c3;
        10'h127: oHanning = 16'h13dc;
        10'h128: oHanning = 16'h13f4;
        10'h129: oHanning = 16'h140c;
        10'h12a: oHanning = 16'h1425;
        10'h12b: oHanning = 16'h143d;
        10'h12c: oHanning = 16'h1455;
        10'h12d: oHanning = 16'h146d;
        10'h12e: oHanning = 16'h1485;
        10'h12f: oHanning = 16'h149d;
        10'h130: oHanning = 16'h14b5;
        10'h131: oHanning = 16'h14cd;
        10'h132: oHanning = 16'h14e5;
        10'h133: oHanning = 16'h14fd;
        10'h134: oHanning = 16'h1515;
        10'h135: oHanning = 16'h152d;
        10'h136: oHanning = 16'h1545;
        10'h137: oHanning = 16'h155c;
        10'h138: oHanning = 16'h1574;
        10'h139: oHanning = 16'h158b;
        10'h13a: oHanning = 16'h15a3;
        10'h13b: oHanning = 16'h15ba;
        10'h13c: oHanning = 16'h15d2;
        10'h13d: oHanning = 16'h15e9;
        10'h13e: oHanning = 16'h1600;
        10'h13f: oHanning = 16'h1618;
        10'h140: oHanning = 16'h162f;
        10'h141: oHanning = 16'h1646;
        10'h142: oHanning = 16'h165d;
        10'h143: oHanning = 16'h1674;
        10'h144: oHanning = 16'h168b;
        10'h145: oHanning = 16'h16a2;
        10'h146: oHanning = 16'h16b9;
        10'h147: oHanning = 16'h16cf;
        10'h148: oHanning = 16'h16e6;
        10'h149: oHanning = 16'h16fd;
        10'h14a: oHanning = 16'h1713;
        10'h14b: oHanning = 16'h172a;
        10'h14c: oHanning = 16'h1740;
        10'h14d: oHanning = 16'h1757;
        10'h14e: oHanning = 16'h176d;
        10'h14f: oHanning = 16'h1783;
        10'h150: oHanning = 16'h1799;
        10'h151: oHanning = 16'h17af;
        10'h152: oHanning = 16'h17c5;
        10'h153: oHanning = 16'h17db;
        10'h154: oHanning = 16'h17f1;
        10'h155: oHanning = 16'h1807;
        10'h156: oHanning = 16'h181c;
        10'h157: oHanning = 16'h1832;
        10'h158: oHanning = 16'h1848;
        10'h159: oHanning = 16'h185d;
        10'h15a: oHanning = 16'h1872;
        10'h15b: oHanning = 16'h1888;
        10'h15c: oHanning = 16'h189d;
        10'h15d: oHanning = 16'h18b2;
        10'h15e: oHanning = 16'h18c7;
        10'h15f: oHanning = 16'h18dc;
        10'h160: oHanning = 16'h18f1;
        10'h161: oHanning = 16'h1906;
        10'h162: oHanning = 16'h191a;
        10'h163: oHanning = 16'h192f;
        10'h164: oHanning = 16'h1943;
        10'h165: oHanning = 16'h1958;
        10'h166: oHanning = 16'h196c;
        10'h167: oHanning = 16'h1980;
        10'h168: oHanning = 16'h1995;
        10'h169: oHanning = 16'h19a9;
        10'h16a: oHanning = 16'h19bd;
        10'h16b: oHanning = 16'h19d0;
        10'h16c: oHanning = 16'h19e4;
        10'h16d: oHanning = 16'h19f8;
        10'h16e: oHanning = 16'h1a0c;
        10'h16f: oHanning = 16'h1a1f;
        10'h170: oHanning = 16'h1a32;
        10'h171: oHanning = 16'h1a46;
        10'h172: oHanning = 16'h1a59;
        10'h173: oHanning = 16'h1a6c;
        10'h174: oHanning = 16'h1a7f;
        10'h175: oHanning = 16'h1a92;
        10'h176: oHanning = 16'h1aa5;
        10'h177: oHanning = 16'h1ab7;
        10'h178: oHanning = 16'h1aca;
        10'h179: oHanning = 16'h1adc;
        10'h17a: oHanning = 16'h1aef;
        10'h17b: oHanning = 16'h1b01;
        10'h17c: oHanning = 16'h1b13;
        10'h17d: oHanning = 16'h1b25;
        10'h17e: oHanning = 16'h1b37;
        10'h17f: oHanning = 16'h1b49;
        10'h180: oHanning = 16'h1b5b;
        10'h181: oHanning = 16'h1b6d;
        10'h182: oHanning = 16'h1b7e;
        10'h183: oHanning = 16'h1b8f;
        10'h184: oHanning = 16'h1ba1;
        10'h185: oHanning = 16'h1bb2;
        10'h186: oHanning = 16'h1bc3;
        10'h187: oHanning = 16'h1bd4;
        10'h188: oHanning = 16'h1be5;
        10'h189: oHanning = 16'h1bf6;
        10'h18a: oHanning = 16'h1c06;
        10'h18b: oHanning = 16'h1c17;
        10'h18c: oHanning = 16'h1c27;
        10'h18d: oHanning = 16'h1c37;
        10'h18e: oHanning = 16'h1c47;
        10'h18f: oHanning = 16'h1c58;
        10'h190: oHanning = 16'h1c67;
        10'h191: oHanning = 16'h1c77;
        10'h192: oHanning = 16'h1c87;
        10'h193: oHanning = 16'h1c96;
        10'h194: oHanning = 16'h1ca6;
        10'h195: oHanning = 16'h1cb5;
        10'h196: oHanning = 16'h1cc4;
        10'h197: oHanning = 16'h1cd3;
        10'h198: oHanning = 16'h1ce2;
        10'h199: oHanning = 16'h1cf1;
        10'h19a: oHanning = 16'h1d00;
        10'h19b: oHanning = 16'h1d0f;
        10'h19c: oHanning = 16'h1d1d;
        10'h19d: oHanning = 16'h1d2b;
        10'h19e: oHanning = 16'h1d39;
        10'h19f: oHanning = 16'h1d48;
        10'h1a0: oHanning = 16'h1d55;
        10'h1a1: oHanning = 16'h1d63;
        10'h1a2: oHanning = 16'h1d71;
        10'h1a3: oHanning = 16'h1d7e;
        10'h1a4: oHanning = 16'h1d8c;
        10'h1a5: oHanning = 16'h1d99;
        10'h1a6: oHanning = 16'h1da6;
        10'h1a7: oHanning = 16'h1db3;
        10'h1a8: oHanning = 16'h1dc0;
        10'h1a9: oHanning = 16'h1dcd;
        10'h1aa: oHanning = 16'h1dda;
        10'h1ab: oHanning = 16'h1de6;
        10'h1ac: oHanning = 16'h1df3;
        10'h1ad: oHanning = 16'h1dff;
        10'h1ae: oHanning = 16'h1e0b;
        10'h1af: oHanning = 16'h1e17;
        10'h1b0: oHanning = 16'h1e23;
        10'h1b1: oHanning = 16'h1e2e;
        10'h1b2: oHanning = 16'h1e3a;
        10'h1b3: oHanning = 16'h1e45;
        10'h1b4: oHanning = 16'h1e51;
        10'h1b5: oHanning = 16'h1e5c;
        10'h1b6: oHanning = 16'h1e67;
        10'h1b7: oHanning = 16'h1e72;
        10'h1b8: oHanning = 16'h1e7c;
        10'h1b9: oHanning = 16'h1e87;
        10'h1ba: oHanning = 16'h1e91;
        10'h1bb: oHanning = 16'h1e9c;
        10'h1bc: oHanning = 16'h1ea6;
        10'h1bd: oHanning = 16'h1eb0;
        10'h1be: oHanning = 16'h1eba;
        10'h1bf: oHanning = 16'h1ec3;
        10'h1c0: oHanning = 16'h1ecd;
        10'h1c1: oHanning = 16'h1ed7;
        10'h1c2: oHanning = 16'h1ee0;
        10'h1c3: oHanning = 16'h1ee9;
        10'h1c4: oHanning = 16'h1ef2;
        10'h1c5: oHanning = 16'h1efb;
        10'h1c6: oHanning = 16'h1f04;
        10'h1c7: oHanning = 16'h1f0c;
        10'h1c8: oHanning = 16'h1f15;
        10'h1c9: oHanning = 16'h1f1d;
        10'h1ca: oHanning = 16'h1f25;
        10'h1cb: oHanning = 16'h1f2d;
        10'h1cc: oHanning = 16'h1f35;
        10'h1cd: oHanning = 16'h1f3d;
        10'h1ce: oHanning = 16'h1f44;
        10'h1cf: oHanning = 16'h1f4c;
        10'h1d0: oHanning = 16'h1f53;
        10'h1d1: oHanning = 16'h1f5a;
        10'h1d2: oHanning = 16'h1f61;
        10'h1d3: oHanning = 16'h1f68;
        10'h1d4: oHanning = 16'h1f6f;
        10'h1d5: oHanning = 16'h1f75;
        10'h1d6: oHanning = 16'h1f7c;
        10'h1d7: oHanning = 16'h1f82;
        10'h1d8: oHanning = 16'h1f88;
        10'h1d9: oHanning = 16'h1f8e;
        10'h1da: oHanning = 16'h1f94;
        10'h1db: oHanning = 16'h1f99;
        10'h1dc: oHanning = 16'h1f9f;
        10'h1dd: oHanning = 16'h1fa4;
        10'h1de: oHanning = 16'h1fa9;
        10'h1df: oHanning = 16'h1fae;
        10'h1e0: oHanning = 16'h1fb3;
        10'h1e1: oHanning = 16'h1fb8;
        10'h1e2: oHanning = 16'h1fbd;
        10'h1e3: oHanning = 16'h1fc1;
        10'h1e4: oHanning = 16'h1fc5;
        10'h1e5: oHanning = 16'h1fca;
        10'h1e6: oHanning = 16'h1fce;
        10'h1e7: oHanning = 16'h1fd1;
        10'h1e8: oHanning = 16'h1fd5;
        10'h1e9: oHanning = 16'h1fd9;
        10'h1ea: oHanning = 16'h1fdc;
        10'h1eb: oHanning = 16'h1fdf;
        10'h1ec: oHanning = 16'h1fe2;
        10'h1ed: oHanning = 16'h1fe5;
        10'h1ee: oHanning = 16'h1fe8;
        10'h1ef: oHanning = 16'h1feb;
        10'h1f0: oHanning = 16'h1fed;
        10'h1f1: oHanning = 16'h1fef;
        10'h1f2: oHanning = 16'h1ff1;
        10'h1f3: oHanning = 16'h1ff3;
        10'h1f4: oHanning = 16'h1ff5;
        10'h1f5: oHanning = 16'h1ff7;
        10'h1f6: oHanning = 16'h1ff9;
        10'h1f7: oHanning = 16'h1ffa;
        10'h1f8: oHanning = 16'h1ffb;
        10'h1f9: oHanning = 16'h1ffc;
        10'h1fa: oHanning = 16'h1ffd;
        10'h1fb: oHanning = 16'h1ffe;
        10'h1fc: oHanning = 16'h1fff;
        10'h1fd: oHanning = 16'h1fff;
        10'h1fe: oHanning = 16'h1fff;
        10'h1ff: oHanning = 16'h1fff;
        10'h200: oHanning = 16'h1fff;
        10'h201: oHanning = 16'h1fff;
        10'h202: oHanning = 16'h1fff;
        10'h203: oHanning = 16'h1fff;
        10'h204: oHanning = 16'h1ffe;
        10'h205: oHanning = 16'h1ffd;
        10'h206: oHanning = 16'h1ffc;
        10'h207: oHanning = 16'h1ffb;
        10'h208: oHanning = 16'h1ffa;
        10'h209: oHanning = 16'h1ff9;
        10'h20a: oHanning = 16'h1ff7;
        10'h20b: oHanning = 16'h1ff5;
        10'h20c: oHanning = 16'h1ff3;
        10'h20d: oHanning = 16'h1ff1;
        10'h20e: oHanning = 16'h1fef;
        10'h20f: oHanning = 16'h1fed;
        10'h210: oHanning = 16'h1feb;
        10'h211: oHanning = 16'h1fe8;
        10'h212: oHanning = 16'h1fe5;
        10'h213: oHanning = 16'h1fe2;
        10'h214: oHanning = 16'h1fdf;
        10'h215: oHanning = 16'h1fdc;
        10'h216: oHanning = 16'h1fd9;
        10'h217: oHanning = 16'h1fd5;
        10'h218: oHanning = 16'h1fd1;
        10'h219: oHanning = 16'h1fce;
        10'h21a: oHanning = 16'h1fca;
        10'h21b: oHanning = 16'h1fc5;
        10'h21c: oHanning = 16'h1fc1;
        10'h21d: oHanning = 16'h1fbd;
        10'h21e: oHanning = 16'h1fb8;
        10'h21f: oHanning = 16'h1fb3;
        10'h220: oHanning = 16'h1fae;
        10'h221: oHanning = 16'h1fa9;
        10'h222: oHanning = 16'h1fa4;
        10'h223: oHanning = 16'h1f9f;
        10'h224: oHanning = 16'h1f99;
        10'h225: oHanning = 16'h1f94;
        10'h226: oHanning = 16'h1f8e;
        10'h227: oHanning = 16'h1f88;
        10'h228: oHanning = 16'h1f82;
        10'h229: oHanning = 16'h1f7c;
        10'h22a: oHanning = 16'h1f75;
        10'h22b: oHanning = 16'h1f6f;
        10'h22c: oHanning = 16'h1f68;
        10'h22d: oHanning = 16'h1f61;
        10'h22e: oHanning = 16'h1f5a;
        10'h22f: oHanning = 16'h1f53;
        10'h230: oHanning = 16'h1f4c;
        10'h231: oHanning = 16'h1f44;
        10'h232: oHanning = 16'h1f3d;
        10'h233: oHanning = 16'h1f35;
        10'h234: oHanning = 16'h1f2d;
        10'h235: oHanning = 16'h1f25;
        10'h236: oHanning = 16'h1f1d;
        10'h237: oHanning = 16'h1f15;
        10'h238: oHanning = 16'h1f0c;
        10'h239: oHanning = 16'h1f04;
        10'h23a: oHanning = 16'h1efb;
        10'h23b: oHanning = 16'h1ef2;
        10'h23c: oHanning = 16'h1ee9;
        10'h23d: oHanning = 16'h1ee0;
        10'h23e: oHanning = 16'h1ed7;
        10'h23f: oHanning = 16'h1ecd;
        10'h240: oHanning = 16'h1ec3;
        10'h241: oHanning = 16'h1eba;
        10'h242: oHanning = 16'h1eb0;
        10'h243: oHanning = 16'h1ea6;
        10'h244: oHanning = 16'h1e9c;
        10'h245: oHanning = 16'h1e91;
        10'h246: oHanning = 16'h1e87;
        10'h247: oHanning = 16'h1e7c;
        10'h248: oHanning = 16'h1e72;
        10'h249: oHanning = 16'h1e67;
        10'h24a: oHanning = 16'h1e5c;
        10'h24b: oHanning = 16'h1e51;
        10'h24c: oHanning = 16'h1e45;
        10'h24d: oHanning = 16'h1e3a;
        10'h24e: oHanning = 16'h1e2e;
        10'h24f: oHanning = 16'h1e23;
        10'h250: oHanning = 16'h1e17;
        10'h251: oHanning = 16'h1e0b;
        10'h252: oHanning = 16'h1dff;
        10'h253: oHanning = 16'h1df3;
        10'h254: oHanning = 16'h1de6;
        10'h255: oHanning = 16'h1dda;
        10'h256: oHanning = 16'h1dcd;
        10'h257: oHanning = 16'h1dc0;
        10'h258: oHanning = 16'h1db3;
        10'h259: oHanning = 16'h1da6;
        10'h25a: oHanning = 16'h1d99;
        10'h25b: oHanning = 16'h1d8c;
        10'h25c: oHanning = 16'h1d7e;
        10'h25d: oHanning = 16'h1d71;
        10'h25e: oHanning = 16'h1d63;
        10'h25f: oHanning = 16'h1d55;
        10'h260: oHanning = 16'h1d48;
        10'h261: oHanning = 16'h1d39;
        10'h262: oHanning = 16'h1d2b;
        10'h263: oHanning = 16'h1d1d;
        10'h264: oHanning = 16'h1d0f;
        10'h265: oHanning = 16'h1d00;
        10'h266: oHanning = 16'h1cf1;
        10'h267: oHanning = 16'h1ce2;
        10'h268: oHanning = 16'h1cd3;
        10'h269: oHanning = 16'h1cc4;
        10'h26a: oHanning = 16'h1cb5;
        10'h26b: oHanning = 16'h1ca6;
        10'h26c: oHanning = 16'h1c96;
        10'h26d: oHanning = 16'h1c87;
        10'h26e: oHanning = 16'h1c77;
        10'h26f: oHanning = 16'h1c67;
        10'h270: oHanning = 16'h1c58;
        10'h271: oHanning = 16'h1c47;
        10'h272: oHanning = 16'h1c37;
        10'h273: oHanning = 16'h1c27;
        10'h274: oHanning = 16'h1c17;
        10'h275: oHanning = 16'h1c06;
        10'h276: oHanning = 16'h1bf6;
        10'h277: oHanning = 16'h1be5;
        10'h278: oHanning = 16'h1bd4;
        10'h279: oHanning = 16'h1bc3;
        10'h27a: oHanning = 16'h1bb2;
        10'h27b: oHanning = 16'h1ba1;
        10'h27c: oHanning = 16'h1b8f;
        10'h27d: oHanning = 16'h1b7e;
        10'h27e: oHanning = 16'h1b6d;
        10'h27f: oHanning = 16'h1b5b;
        10'h280: oHanning = 16'h1b49;
        10'h281: oHanning = 16'h1b37;
        10'h282: oHanning = 16'h1b25;
        10'h283: oHanning = 16'h1b13;
        10'h284: oHanning = 16'h1b01;
        10'h285: oHanning = 16'h1aef;
        10'h286: oHanning = 16'h1adc;
        10'h287: oHanning = 16'h1aca;
        10'h288: oHanning = 16'h1ab7;
        10'h289: oHanning = 16'h1aa5;
        10'h28a: oHanning = 16'h1a92;
        10'h28b: oHanning = 16'h1a7f;
        10'h28c: oHanning = 16'h1a6c;
        10'h28d: oHanning = 16'h1a59;
        10'h28e: oHanning = 16'h1a46;
        10'h28f: oHanning = 16'h1a32;
        10'h290: oHanning = 16'h1a1f;
        10'h291: oHanning = 16'h1a0c;
        10'h292: oHanning = 16'h19f8;
        10'h293: oHanning = 16'h19e4;
        10'h294: oHanning = 16'h19d0;
        10'h295: oHanning = 16'h19bd;
        10'h296: oHanning = 16'h19a9;
        10'h297: oHanning = 16'h1995;
        10'h298: oHanning = 16'h1980;
        10'h299: oHanning = 16'h196c;
        10'h29a: oHanning = 16'h1958;
        10'h29b: oHanning = 16'h1943;
        10'h29c: oHanning = 16'h192f;
        10'h29d: oHanning = 16'h191a;
        10'h29e: oHanning = 16'h1906;
        10'h29f: oHanning = 16'h18f1;
        10'h2a0: oHanning = 16'h18dc;
        10'h2a1: oHanning = 16'h18c7;
        10'h2a2: oHanning = 16'h18b2;
        10'h2a3: oHanning = 16'h189d;
        10'h2a4: oHanning = 16'h1888;
        10'h2a5: oHanning = 16'h1872;
        10'h2a6: oHanning = 16'h185d;
        10'h2a7: oHanning = 16'h1848;
        10'h2a8: oHanning = 16'h1832;
        10'h2a9: oHanning = 16'h181c;
        10'h2aa: oHanning = 16'h1807;
        10'h2ab: oHanning = 16'h17f1;
        10'h2ac: oHanning = 16'h17db;
        10'h2ad: oHanning = 16'h17c5;
        10'h2ae: oHanning = 16'h17af;
        10'h2af: oHanning = 16'h1799;
        10'h2b0: oHanning = 16'h1783;
        10'h2b1: oHanning = 16'h176d;
        10'h2b2: oHanning = 16'h1757;
        10'h2b3: oHanning = 16'h1740;
        10'h2b4: oHanning = 16'h172a;
        10'h2b5: oHanning = 16'h1713;
        10'h2b6: oHanning = 16'h16fd;
        10'h2b7: oHanning = 16'h16e6;
        10'h2b8: oHanning = 16'h16cf;
        10'h2b9: oHanning = 16'h16b9;
        10'h2ba: oHanning = 16'h16a2;
        10'h2bb: oHanning = 16'h168b;
        10'h2bc: oHanning = 16'h1674;
        10'h2bd: oHanning = 16'h165d;
        10'h2be: oHanning = 16'h1646;
        10'h2bf: oHanning = 16'h162f;
        10'h2c0: oHanning = 16'h1618;
        10'h2c1: oHanning = 16'h1600;
        10'h2c2: oHanning = 16'h15e9;
        10'h2c3: oHanning = 16'h15d2;
        10'h2c4: oHanning = 16'h15ba;
        10'h2c5: oHanning = 16'h15a3;
        10'h2c6: oHanning = 16'h158b;
        10'h2c7: oHanning = 16'h1574;
        10'h2c8: oHanning = 16'h155c;
        10'h2c9: oHanning = 16'h1545;
        10'h2ca: oHanning = 16'h152d;
        10'h2cb: oHanning = 16'h1515;
        10'h2cc: oHanning = 16'h14fd;
        10'h2cd: oHanning = 16'h14e5;
        10'h2ce: oHanning = 16'h14cd;
        10'h2cf: oHanning = 16'h14b5;
        10'h2d0: oHanning = 16'h149d;
        10'h2d1: oHanning = 16'h1485;
        10'h2d2: oHanning = 16'h146d;
        10'h2d3: oHanning = 16'h1455;
        10'h2d4: oHanning = 16'h143d;
        10'h2d5: oHanning = 16'h1425;
        10'h2d6: oHanning = 16'h140c;
        10'h2d7: oHanning = 16'h13f4;
        10'h2d8: oHanning = 16'h13dc;
        10'h2d9: oHanning = 16'h13c3;
        10'h2da: oHanning = 16'h13ab;
        10'h2db: oHanning = 16'h1392;
        10'h2dc: oHanning = 16'h137a;
        10'h2dd: oHanning = 16'h1361;
        10'h2de: oHanning = 16'h1349;
        10'h2df: oHanning = 16'h1330;
        10'h2e0: oHanning = 16'h1318;
        10'h2e1: oHanning = 16'h12ff;
        10'h2e2: oHanning = 16'h12e6;
        10'h2e3: oHanning = 16'h12ce;
        10'h2e4: oHanning = 16'h12b5;
        10'h2e5: oHanning = 16'h129c;
        10'h2e6: oHanning = 16'h1283;
        10'h2e7: oHanning = 16'h126b;
        10'h2e8: oHanning = 16'h1252;
        10'h2e9: oHanning = 16'h1239;
        10'h2ea: oHanning = 16'h1220;
        10'h2eb: oHanning = 16'h1207;
        10'h2ec: oHanning = 16'h11ee;
        10'h2ed: oHanning = 16'h11d5;
        10'h2ee: oHanning = 16'h11bc;
        10'h2ef: oHanning = 16'h11a3;
        10'h2f0: oHanning = 16'h118a;
        10'h2f1: oHanning = 16'h1171;
        10'h2f2: oHanning = 16'h1158;
        10'h2f3: oHanning = 16'h113f;
        10'h2f4: oHanning = 16'h1126;
        10'h2f5: oHanning = 16'h110d;
        10'h2f6: oHanning = 16'h10f4;
        10'h2f7: oHanning = 16'h10db;
        10'h2f8: oHanning = 16'h10c2;
        10'h2f9: oHanning = 16'h10a9;
        10'h2fa: oHanning = 16'h1090;
        10'h2fb: oHanning = 16'h1077;
        10'h2fc: oHanning = 16'h105e;
        10'h2fd: oHanning = 16'h1045;
        10'h2fe: oHanning = 16'h102b;
        10'h2ff: oHanning = 16'h1012;
        10'h300: oHanning = 16'hff9;
        10'h301: oHanning = 16'hfe0;
        10'h302: oHanning = 16'hfc7;
        10'h303: oHanning = 16'hfae;
        10'h304: oHanning = 16'hf95;
        10'h305: oHanning = 16'hf7c;
        10'h306: oHanning = 16'hf63;
        10'h307: oHanning = 16'hf4a;
        10'h308: oHanning = 16'hf30;
        10'h309: oHanning = 16'hf17;
        10'h30a: oHanning = 16'hefe;
        10'h30b: oHanning = 16'hee5;
        10'h30c: oHanning = 16'hecc;
        10'h30d: oHanning = 16'heb3;
        10'h30e: oHanning = 16'he9a;
        10'h30f: oHanning = 16'he81;
        10'h310: oHanning = 16'he68;
        10'h311: oHanning = 16'he4f;
        10'h312: oHanning = 16'he36;
        10'h313: oHanning = 16'he1d;
        10'h314: oHanning = 16'he04;
        10'h315: oHanning = 16'hdeb;
        10'h316: oHanning = 16'hdd3;
        10'h317: oHanning = 16'hdba;
        10'h318: oHanning = 16'hda1;
        10'h319: oHanning = 16'hd88;
        10'h31a: oHanning = 16'hd6f;
        10'h31b: oHanning = 16'hd56;
        10'h31c: oHanning = 16'hd3e;
        10'h31d: oHanning = 16'hd25;
        10'h31e: oHanning = 16'hd0c;
        10'h31f: oHanning = 16'hcf4;
        10'h320: oHanning = 16'hcdb;
        10'h321: oHanning = 16'hcc2;
        10'h322: oHanning = 16'hcaa;
        10'h323: oHanning = 16'hc91;
        10'h324: oHanning = 16'hc79;
        10'h325: oHanning = 16'hc60;
        10'h326: oHanning = 16'hc48;
        10'h327: oHanning = 16'hc2f;
        10'h328: oHanning = 16'hc17;
        10'h329: oHanning = 16'hbff;
        10'h32a: oHanning = 16'hbe6;
        10'h32b: oHanning = 16'hbce;
        10'h32c: oHanning = 16'hbb6;
        10'h32d: oHanning = 16'hb9e;
        10'h32e: oHanning = 16'hb86;
        10'h32f: oHanning = 16'hb6e;
        10'h330: oHanning = 16'hb56;
        10'h331: oHanning = 16'hb3e;
        10'h332: oHanning = 16'hb26;
        10'h333: oHanning = 16'hb0e;
        10'h334: oHanning = 16'haf6;
        10'h335: oHanning = 16'hade;
        10'h336: oHanning = 16'hac6;
        10'h337: oHanning = 16'haaf;
        10'h338: oHanning = 16'ha97;
        10'h339: oHanning = 16'ha7f;
        10'h33a: oHanning = 16'ha68;
        10'h33b: oHanning = 16'ha50;
        10'h33c: oHanning = 16'ha39;
        10'h33d: oHanning = 16'ha21;
        10'h33e: oHanning = 16'ha0a;
        10'h33f: oHanning = 16'h9f3;
        10'h340: oHanning = 16'h9dc;
        10'h341: oHanning = 16'h9c5;
        10'h342: oHanning = 16'h9ad;
        10'h343: oHanning = 16'h996;
        10'h344: oHanning = 16'h97f;
        10'h345: oHanning = 16'h969;
        10'h346: oHanning = 16'h952;
        10'h347: oHanning = 16'h93b;
        10'h348: oHanning = 16'h924;
        10'h349: oHanning = 16'h90e;
        10'h34a: oHanning = 16'h8f7;
        10'h34b: oHanning = 16'h8e0;
        10'h34c: oHanning = 16'h8ca;
        10'h34d: oHanning = 16'h8b4;
        10'h34e: oHanning = 16'h89d;
        10'h34f: oHanning = 16'h887;
        10'h350: oHanning = 16'h871;
        10'h351: oHanning = 16'h85b;
        10'h352: oHanning = 16'h845;
        10'h353: oHanning = 16'h82f;
        10'h354: oHanning = 16'h819;
        10'h355: oHanning = 16'h803;
        10'h356: oHanning = 16'h7ed;
        10'h357: oHanning = 16'h7d8;
        10'h358: oHanning = 16'h7c2;
        10'h359: oHanning = 16'h7ad;
        10'h35a: oHanning = 16'h797;
        10'h35b: oHanning = 16'h782;
        10'h35c: oHanning = 16'h76d;
        10'h35d: oHanning = 16'h758;
        10'h35e: oHanning = 16'h743;
        10'h35f: oHanning = 16'h72e;
        10'h360: oHanning = 16'h719;
        10'h361: oHanning = 16'h704;
        10'h362: oHanning = 16'h6ef;
        10'h363: oHanning = 16'h6da;
        10'h364: oHanning = 16'h6c6;
        10'h365: oHanning = 16'h6b1;
        10'h366: oHanning = 16'h69d;
        10'h367: oHanning = 16'h689;
        10'h368: oHanning = 16'h675;
        10'h369: oHanning = 16'h660;
        10'h36a: oHanning = 16'h64c;
        10'h36b: oHanning = 16'h638;
        10'h36c: oHanning = 16'h625;
        10'h36d: oHanning = 16'h611;
        10'h36e: oHanning = 16'h5fd;
        10'h36f: oHanning = 16'h5ea;
        10'h370: oHanning = 16'h5d6;
        10'h371: oHanning = 16'h5c3;
        10'h372: oHanning = 16'h5b0;
        10'h373: oHanning = 16'h59d;
        10'h374: oHanning = 16'h58a;
        10'h375: oHanning = 16'h577;
        10'h376: oHanning = 16'h564;
        10'h377: oHanning = 16'h551;
        10'h378: oHanning = 16'h53e;
        10'h379: oHanning = 16'h52c;
        10'h37a: oHanning = 16'h519;
        10'h37b: oHanning = 16'h507;
        10'h37c: oHanning = 16'h4f5;
        10'h37d: oHanning = 16'h4e3;
        10'h37e: oHanning = 16'h4d1;
        10'h37f: oHanning = 16'h4bf;
        10'h380: oHanning = 16'h4ad;
        10'h381: oHanning = 16'h49b;
        10'h382: oHanning = 16'h48a;
        10'h383: oHanning = 16'h478;
        10'h384: oHanning = 16'h467;
        10'h385: oHanning = 16'h456;
        10'h386: oHanning = 16'h445;
        10'h387: oHanning = 16'h433;
        10'h388: oHanning = 16'h423;
        10'h389: oHanning = 16'h412;
        10'h38a: oHanning = 16'h401;
        10'h38b: oHanning = 16'h3f1;
        10'h38c: oHanning = 16'h3e0;
        10'h38d: oHanning = 16'h3d0;
        10'h38e: oHanning = 16'h3c0;
        10'h38f: oHanning = 16'h3af;
        10'h390: oHanning = 16'h3a0;
        10'h391: oHanning = 16'h390;
        10'h392: oHanning = 16'h380;
        10'h393: oHanning = 16'h370;
        10'h394: oHanning = 16'h361;
        10'h395: oHanning = 16'h351;
        10'h396: oHanning = 16'h342;
        10'h397: oHanning = 16'h333;
        10'h398: oHanning = 16'h324;
        10'h399: oHanning = 16'h315;
        10'h39a: oHanning = 16'h306;
        10'h39b: oHanning = 16'h2f8;
        10'h39c: oHanning = 16'h2e9;
        10'h39d: oHanning = 16'h2db;
        10'h39e: oHanning = 16'h2cd;
        10'h39f: oHanning = 16'h2be;
        10'h3a0: oHanning = 16'h2b0;
        10'h3a1: oHanning = 16'h2a3;
        10'h3a2: oHanning = 16'h295;
        10'h3a3: oHanning = 16'h287;
        10'h3a4: oHanning = 16'h27a;
        10'h3a5: oHanning = 16'h26c;
        10'h3a6: oHanning = 16'h25f;
        10'h3a7: oHanning = 16'h252;
        10'h3a8: oHanning = 16'h245;
        10'h3a9: oHanning = 16'h238;
        10'h3aa: oHanning = 16'h22c;
        10'h3ab: oHanning = 16'h21f;
        10'h3ac: oHanning = 16'h213;
        10'h3ad: oHanning = 16'h206;
        10'h3ae: oHanning = 16'h1fa;
        10'h3af: oHanning = 16'h1ee;
        10'h3b0: oHanning = 16'h1e2;
        10'h3b1: oHanning = 16'h1d6;
        10'h3b2: oHanning = 16'h1cb;
        10'h3b3: oHanning = 16'h1bf;
        10'h3b4: oHanning = 16'h1b4;
        10'h3b5: oHanning = 16'h1a9;
        10'h3b6: oHanning = 16'h19e;
        10'h3b7: oHanning = 16'h193;
        10'h3b8: oHanning = 16'h188;
        10'h3b9: oHanning = 16'h17d;
        10'h3ba: oHanning = 16'h173;
        10'h3bb: oHanning = 16'h168;
        10'h3bc: oHanning = 16'h15e;
        10'h3bd: oHanning = 16'h154;
        10'h3be: oHanning = 16'h14a;
        10'h3bf: oHanning = 16'h140;
        10'h3c0: oHanning = 16'h137;
        10'h3c1: oHanning = 16'h12d;
        10'h3c2: oHanning = 16'h124;
        10'h3c3: oHanning = 16'h11b;
        10'h3c4: oHanning = 16'h111;
        10'h3c5: oHanning = 16'h108;
        10'h3c6: oHanning = 16'h100;
        10'h3c7: oHanning = 16'h0f7;
        10'h3c8: oHanning = 16'h0ee;
        10'h3c9: oHanning = 16'h0e6;
        10'h3ca: oHanning = 16'h0de;
        10'h3cb: oHanning = 16'h0d6;
        10'h3cc: oHanning = 16'h0ce;
        10'h3cd: oHanning = 16'h0c6;
        10'h3ce: oHanning = 16'h0be;
        10'h3cf: oHanning = 16'h0b7;
        10'h3d0: oHanning = 16'h0b0;
        10'h3d1: oHanning = 16'h0a8;
        10'h3d2: oHanning = 16'h0a1;
        10'h3d3: oHanning = 16'h09a;
        10'h3d4: oHanning = 16'h094;
        10'h3d5: oHanning = 16'h08d;
        10'h3d6: oHanning = 16'h087;
        10'h3d7: oHanning = 16'h080;
        10'h3d8: oHanning = 16'h07a;
        10'h3d9: oHanning = 16'h074;
        10'h3da: oHanning = 16'h06e;
        10'h3db: oHanning = 16'h068;
        10'h3dc: oHanning = 16'h063;
        10'h3dd: oHanning = 16'h05d;
        10'h3de: oHanning = 16'h058;
        10'h3df: oHanning = 16'h053;
        10'h3e0: oHanning = 16'h04e;
        10'h3e1: oHanning = 16'h049;
        10'h3e2: oHanning = 16'h045;
        10'h3e3: oHanning = 16'h040;
        10'h3e4: oHanning = 16'h03c;
        10'h3e5: oHanning = 16'h037;
        10'h3e6: oHanning = 16'h033;
        10'h3e7: oHanning = 16'h030;
        10'h3e8: oHanning = 16'h02c;
        10'h3e9: oHanning = 16'h028;
        10'h3ea: oHanning = 16'h025;
        10'h3eb: oHanning = 16'h021;
        10'h3ec: oHanning = 16'h01e;
        10'h3ed: oHanning = 16'h01b;
        10'h3ee: oHanning = 16'h018;
        10'h3ef: oHanning = 16'h016;
        10'h3f0: oHanning = 16'h013;
        10'h3f1: oHanning = 16'h011;
        10'h3f2: oHanning = 16'h00f;
        10'h3f3: oHanning = 16'h00c;
        10'h3f4: oHanning = 16'h00b;
        10'h3f5: oHanning = 16'h009;
        10'h3f6: oHanning = 16'h007;
        10'h3f7: oHanning = 16'h006;
        10'h3f8: oHanning = 16'h004;
        10'h3f9: oHanning = 16'h003;
        10'h3fa: oHanning = 16'h002;
        10'h3fb: oHanning = 16'h001;
        10'h3fc: oHanning = 16'h001;
        10'h3fd: oHanning = 16'h000;
        10'h3fe: oHanning = 16'h000;
        10'h3ff: oHanning = 16'h000;
    endcase
end

endmodule